----------------------------------------------------------------------------------
-- Company: Vaga SA
-- Engineer: Mamoyano
-- 
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

entity rom_meta is
	generic (
		ADDRESS_WIDE : integer := 8;
		DATA_WIDE : integer := 2
	);
	port(
		clk1: in std_logic;
		we1 : in std_logic;
		input1 : in std_logic_vector(DATA_WIDE - 1 downto 0); --(DATA_WIDE - 1 downto 0)
		addr1 : in std_logic_vector(ADDRESS_WIDE - 1 downto 0);
		salida1 : out std_logic_vector(DATA_WIDE - 1 downto 0)
	);
end rom_meta;

architecture Behavioral of rom_meta is
	
	type TMemory is array (0 to 2** ADDRESS_WIDE - 1) of std_logic_vector(DATA_WIDE - 1 downto 0);

	shared variable memory : TMemory := 
	( 
		"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
		"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
		"00","00","00","00","10","10","10","10","10","10","10","10","00","00","00","00",
		"00","00","00","00","00","10","10","10","10","10","10","00","00","00","00","00",
		"00","00","10","10","00","10","10","10","10","10","10","00","10","10","00","00",
		"00","00","10","00","10","10","10","10","10","10","10","10","00","10","00","00",
		"00","00","10","00","00","10","10","10","10","10","10","00","00","10","00","00",
		"00","00","10","00","00","10","10","10","10","10","10","00","00","10","00","00",
		"00","00","00","10","00","10","10","10","10","10","10","00","10","00","00","00",
		"00","00","00","00","10","10","10","10","10","10","10","10","00","00","00","00",
		"00","00","00","00","00","10","10","10","10","10","10","00","00","00","00","00",
		"00","00","00","00","00","10","10","10","10","10","10","00","00","00","00","00",
		"00","00","00","00","00","00","10","10","10","10","00","00","00","00","00","00",
		"00","00","00","00","10","10","10","10","10","10","10","10","00","00","00","00",
		"00","00","00","10","10","10","10","10","10","10","10","10","10","00","00","00",
		"00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00"
		
	);

begin

	process (clk1) -- Process de la ROM
	begin

		if clk1'event and clk1 = '1' then
			if we1 = '1' then
				memory(conv_integer(addr1)) := input1;
			end if;
			salida1 <= memory(conv_integer(addr1));
		end if;
	end process;

											
end Behavioral;